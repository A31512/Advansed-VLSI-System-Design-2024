`define R_TYPE    7'b0110011
`define I_TYPE    7'b0010011
`define LOAD      7'b0000011
`define JALR      7'b1100111
`define STORE     7'b0100011
`define B_TYPE    7'b1100011
`define AUPIC     7'b0010111
`define LUI       7'b0110111
`define JAL       7'b1101111
`define FSW       7'b0100111
`define FLW       7'b0000111
`define F_TYPE    7'b1010011 //83
`define CSR_TYPE  7'b1110011 

`define ADD    5'b00000
`define SUB    5'b00010
`define SLL    5'b00100
`define SLT    5'b01000
`define SLTU   5'b01100
`define XOR    5'b10000
`define SRL    5'b10100
`define SRA    5'b10110
`define OR     5'b11000
`define AND    5'b11100
`define MUL    5'b00001
`define MULH   5'b00101
`define MULHU  5'b01001
`define MULHSU 5'b01101
`define FADD   5'b10001 //17
`define FSUB   5'b10101 //21

